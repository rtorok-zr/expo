// Copyright zeroRISC Inc.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

class clk_rst_agent_cfg extends dv_base_agent_cfg;


  `uvm_object_utils_begin(clk_rst_agent_cfg)
  `uvm_object_utils_end

  `uvm_object_new

endclass
